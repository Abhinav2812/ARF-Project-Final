library ieee;
use ieee.std_logic_1164.all;
entity demux1to4 is port(
	S0,S1,S2,S3: OUT STD_LOGIC_VECTOR(15 downto 0);
	sel: IN STD_LOGIC_VECTOR(1 downto 0);
	I: IN STD_LOGIC_VECTOR(15 downto 0)
);
end entity;
architecture behavioral of demux1to4 is
begin
process(I,sel)
begin
	S0 <= x"0000";
	S1 <= x"0000";
	S2 <= x"0000";
	S3 <= x"0000";
	case sel is
	when "00" => S0 <= I;
   when "01" => S1 <= I;
	when "10" => S2 <= I;
   when "11" => S3 <= I;
	end case;
end process;
end architecture;