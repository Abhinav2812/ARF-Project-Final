library verilog;
use verilog.vl_types.all;
entity add_vlg_sample_tst is
    port(
        A               : in     vl_logic_vector(15 downto 0);
        B               : in     vl_logic_vector(15 downto 0);
        en              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end add_vlg_sample_tst;
