library verilog;
use verilog.vl_types.all;
entity demux1to16_vlg_vec_tst is
end demux1to16_vlg_vec_tst;
